<?xml version="1.0" encoding="UTF-8"?>
<svg width="1280" height="320" viewBox="0 0 1280 320" role="img" xmlns="http://www.w3.org/2000/svg" aria-labelledby="title desc">
  <title id="title">Hanu Dixit — Quantum-safe SMPC • Cybersecurity • PM</title>
  <desc id="desc">A clean, geometric banner with subtle quantum motif and high contrast text.</desc>
  <defs>
    <linearGradient id="g" x1="0" y1="0" x2="1" y2="1">
      <stop offset="0%" stop-color="#0f172a"/>
      <stop offset="100%" stop-color="#111827"/>
    </linearGradient>
    <pattern id="qp" x="0" y="0" width="40" height="40" patternUnits="userSpaceOnUse">
      <circle cx="20" cy="20" r="1.5" fill="#475569" opacity="0.35"/>
      <path d="M20 0 L20 40 M0 20 L40 20" stroke="#334155" stroke-width="0.25" opacity="0.25"/>
    </pattern>
  </defs>

  <rect width="1280" height="320" fill="url(#g)"/>
  <rect width="1280" height="320" fill="url(#qp)" opacity="0.35"/>

  <g opacity="0.25">
    <g transform="translate(980,70)">
      <polygon points="0,0 80,0 120,35 40,35" fill="#22d3ee" opacity="0.15"/>
      <polygon points="40,35 120,35 160,70 80,70" fill="#a78bfa" opacity="0.15"/>
      <polygon points="80,70 160,70 200,105 120,105" fill="#34d399" opacity="0.15"/>
      <circle cx="0" cy="0" r="3" fill="#22d3ee"/>
      <circle cx="80" cy="0" r="3" fill="#22d3ee"/>
      <circle cx="120" cy="35" r="3" fill="#a78bfa"/>
      <circle cx="40" cy="35" r="3" fill="#a78bfa"/>
      <circle cx="80" cy="70" r="3" fill="#34d399"/>
      <circle cx="160" cy="70" r="3" fill="#34d399"/>
      <circle cx="200" cy="105" r="3" fill="#34d399"/>
      <circle cx="120" cy="105" r="3" fill="#34d399"/>
      <path d="M0 0 L80 0 L120 35 L40 35 Z M40 35 L120 35 L160 70 L80 70 Z M80 70 L160 70 L200 105 L120 105 Z"
            fill="none" stroke="#cbd5e1" stroke-width="0.6" opacity="0.35"/>
    </g>
  </g>

  <g transform="translate(64,180)">
    <text x="0" y="0" font-family="system-ui,-apple-system,BlinkMacSystemFont,Segoe UI,Roboto,Ubuntu,'Helvetica Neue',Arial" font-size="40" fill="#e5e7eb" font-weight="700">
      Hanu Dixit — Quantum-safe SMPC • Cybersecurity • PM
    </text>
    <text x="0" y="38" font-family="system-ui,-apple-system,BlinkMacSystemFont,Segoe UI,Roboto,Ubuntu,'Helvetica Neue',Arial" font-size="18" fill="#94a3b8">
      Research → Product • PSI • Secure Aggregation • NIST 800-171 nuance
    </text>
  </g>

  <rect x="64" y="208" width="360" height="4" fill="#22d3ee" rx="2"/>
</svg>
